
  

end;

